module alu (
    input  logic [3:0] opcode,
    input  logic [7:0] a, b,
    output logic [15:0] result
);

// Your code here




endmodule


